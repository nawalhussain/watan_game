2
0 0 0 0 0 g c 2 1 
0 0 0 0 0 g c 
0 0 0 0 0 g c 
0 0 0 0 0 g c 
3 8 0 8 4 9 3 4 1 9 3 10 2 4 0 5 0 6 1 6 0 3 5 7 4 11 2 3 2 2 2 11 4 12 1 10 1 5
